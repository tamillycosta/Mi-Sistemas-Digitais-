module hex_to_7segment (
	input clk,
    input  wire [3:0] hex_in,       // Entrada de 4 bits (0 a F)
    output reg  [6:0] seg_out       // Saída para display de 7 segmentos (a-g)
);

//      7 segmentos: seg_out = {a, b, c, d, e, f, g}
// Segmentos ativos em nível baixo (0 = ligado, 1 = desligado)
always @(posedge clk) begin
    case (hex_in)
        4'h0: seg_out = !7'b0000001; // 0
        4'h1: seg_out = !7'b1001111; // 1
        4'h2: seg_out = !7'b0010010; // 2
        4'h3: seg_out = !7'b0000110; // 3
        4'h4: seg_out = !7'b1001100; // 4
        4'h5: seg_out = !7'b0100100; // 5
        4'h6: seg_out = !7'b0100000; // 6
        4'h7: seg_out = !7'b0001111; // 7
        4'h8: seg_out = !7'b0000000; // 8
        4'h9: seg_out = !7'b0000100; // 9
        4'hA: seg_out = !7'b0001000; // A
        4'hB: seg_out = !7'b1100000; // B
        4'hC: seg_out = !7'b0110001; // C
        4'hD: seg_out = !7'b1000010; // D
        4'hE: seg_out = !7'b0110000; // E
        4'hF: seg_out = !7'b0111000; // F
        default: seg_out = !7'b1111111; // Tudo desligado
    endcase
end

endmodule
